module R_subs #(
parameter DW = 16,
parameter DW_2 = 8

) (
input logic [DW_2-1:0] R,
input logic [DW_2-1:0] Q,
output A

);

endmodule